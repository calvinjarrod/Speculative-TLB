`default_nettype wire
module spec_tlb_tb();

// TB TO TLB PORTS
reg TRANS_RQST;
reg SPEC_TLB_RQST;
reg[7:0] VIRT_ADDR_LOOKUP;
wire SPEC_HIT;
wire TLB_HIT;
wire[7:0] PHY_ADDR_TRANS;
wire DONE_TRANS;
reg clk;

// TB TO 8B PT PORTS
reg PT_8B_INSERT_RQST;
reg [4:0] PT_8B_INSERT_INDX;
reg [9:0] PT_8B_INSERT_ENTRY;

// TB TO 32B PT PORTS
reg PT_32B_INSERT_RQST;
reg [3:0] PT_32B_INSERT_INDX;
reg [5:0] PT_32B_INSERT_ENTRY;

// 8B TO TLB INTERCONNECTS
wire LOOKUP_RQST_8B;
wire [4:0] LOOKUP_ADDR_8B;
wire LOOKUP_COMPLETE_8B;
wire [9:0] LOOKUP_RETURN_8B;

// 32B TO TLB INTERCONNECTS
wire LOOKUP_RQST_32B;
wire [2:0] LOOKUP_ADDR_32B;
wire LOOKUP_COMPLETE_32B;
wire [5:0] LOOKUP_RETURN_32B;

SPECLATIVE_TLB SPEC_TLB(
	.SPEC_TLB_RQST(SPEC_TLB_RQST),
	.TRANS_RQST(TRANS_RQST),
	.VIRT_ADDR_LOOKUP(VIRT_ADDR_LOOKUP),
	.SPEC_HIT(SPEC_HIT),
	.TLB_HIT(TLB_HIT),
	.PHY_ADDR_TRANS(PHY_ADDR_TRANS),
	.DONE_TRANS(DONE_TRANS),
	.clk(clk),
	.PAGE_8B_RQST(LOOKUP_RQST_8B),
	.PAGE_8B_LOOKUP(LOOKUP_ADDR_8B),
	.PAGE_8B_RECV(LOOKUP_RETURN_8B),
	.PAGE_8B_COMPLETE(LOOKUP_COMPLETE_8B), 
	.PAGE_32B_RQST(LOOKUP_RQST_32B),
	.PAGE_32B_LOOKUP(LOOKUP_ADDR_32B),
	.PAGE_32B_RECV(LOOKUP_RETURN_32B),
	.PAGE_32B_COMPLETE(LOOKUP_COMPLETE_32B)
);

PAGE_TABLE_32B PT_32B (
	.LOOKUP_RQST(LOOKUP_RQST_32B),
	.LOOKUP_ADDR(LOOKUP_ADDR_32B),
	.LOOKUP_COMPLETE(LOOKUP_COMPLETE_32B),
	.LOOKUP_RETURN(LOOKUP_RETURN_32B),
	.PT_INSERT_RQST(PT_32B_INSERT_RQST),
	.PT_INSERT_INDX(PT_32B_INSERT_INDX),
	.PT_INSERT_ENTRY(PT_32B_INSERT_ENTRY),
	.clk(clk)
);

PAGE_TABLE_8B PT_8B (
	.LOOKUP_RQST(LOOKUP_RQST_8B),
	.LOOKUP_ADDR(LOOKUP_ADDR_8B),
	.LOOKUP_COMPLETE(LOOKUP_COMPLETE_8B),
	.LOOKUP_RETURN(LOOKUP_RETURN_8B),
	.PT_INSERT_RQST(PT_8B_INSERT_RQST),
	.PT_INSERT_INDX(PT_8B_INSERT_INDX),
	.PT_INSERT_ENTRY(PT_8B_INSERT_ENTRY),
	.clk(clk)
);


endmodule
